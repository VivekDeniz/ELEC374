module Not_32(
	input wire [31:0] Ra,
	output wire [31:0] Rz
	);
	//Assign Rz the complement of Ra
	assign Rz = ~Ra ;
	
	
	
endmodule 
