`timescale 1ns/10ps
//OR
module datapath_not_tb;
    reg PCout, ZHighout, Zlowout, Hiout, Loout, InPortout, Cout, MDRout, R2out, R4out;
    reg MARin, PCin, MDRin, IRin, Yin, read, IncPC;
    reg [4:0] opCode;
    reg R5in, R2in, R4in, HIin, LOin, ZHighin, Cin, Zlowin, Clock, Clear;
    reg [31:0] Mdatain;
	 reg branch_flag;
    wire [31:0] reg1out;
    parameter Default = 4'b0000, Reg_load1a = 4'b0001, Reg_load1b = 4'b0010, Reg_load2a = 4'b0011,
             Reg_load2b = 4'b0100, Reg_load3a = 4'b0101, Reg_load3b = 4'b0110, T0 = 4'b0111,
             T1 = 4'b1000, T2 = 4'b1001, T3 = 4'b1010, T4 = 4'b1011, T5 = 4'b1100;
    reg [3:0] Present_state = Default;

    datapath DUT(
        .PCout(PCout), .ZHighout(ZHighout), .Zlowout(Zlowout), .HIout(Hiout), .LOout(Loout), .InPortout(InPortout), .Cout(Cout), .MDRout(MDRout), .R2out(R2out), .R4out(R4out),
        .MARin(MARin), .PCin(PCin), .MDRin(MDRin), .IRin(IRin), .Yin(Yin),
        .IncPC(IncPC), .Read(read), .operation(opCode), .R5in(R5in), .R2in(R2in), .R4in(R4in),
        .clk(Clock), .Mdatain(Mdatain), .clr(Clear), .HIin(HIin), .LOin(LOin), .ZHIin(ZHighin), .ZLOin(ZLOin), .Cin(Cin), .branch_flag(branch_flag), .reg1out(reg1out)
    );

    // Clock generation
    initial begin
        Clear = 0;
        Clock = 0;
        forever #10 Clock = ~Clock; // Toggle clock every 10 time units
    end

    // FSM definition
    always @(posedge Clock) begin
        case (Present_state)
            Default: #40 Present_state = Reg_load1a;
            Reg_load1a: #40 Present_state = Reg_load1b;
            Reg_load1b: #40 Present_state = Reg_load2a;
            Reg_load2a: #40 Present_state = Reg_load2b;
            Reg_load2b: #40 Present_state = Reg_load3a;
            Reg_load3a: #40 Present_state = Reg_load3b;
            Reg_load3b: #40 Present_state = T0;
            T0: #40 Present_state = T1;
            T1: #40 Present_state = T2;
            T2: #40 Present_state = T3;
            T3: #40 Present_state = T4;
            T4: #40 Present_state = T5;
            T5: #40 Present_state = Default; // Reset to default state after T5
        endcase
    end

    // FSM state behavior
    always @(Present_state) begin
        case (Present_state)
            Default: begin
                // Initialize signals
                {PCout, Zlowout, ZHighout, MDRout, R2out, R4out, MARin, Zlowin, PCin, MDRin, IRin, Yin, IncPC, read, branch_flag, Hiout, Loout, InPortout, Cout, R5in, R2in, R4in, Mdatain} = 0;
                opCode = 5'b10010; 
            end
            Reg_load1a: begin
                Mdatain <= 32'h00000012;
                read = 0; MDRin = 0;
                #10; read = 1; MDRin = 1;
                #15; read = 0; MDRin = 0;
            end
            Reg_load1b: begin
                #10; MDRout = 1; R2in = 1;
                #15; MDRout = 0; R2in = 0;
            end
            Reg_load2a: begin
                Mdatain <= 32'h00000014;
                #10; read = 1; MDRin = 1;
                #15; read = 0; MDRin = 0;
            end
            Reg_load2b: begin
                #10; MDRout = 1; R4in = 1;
                #15; MDRout = 0; R4in = 0;
            end
            Reg_load3a: begin
                Mdatain <= 32'h00000018;
                #10; read = 1; MDRin = 1;
                #15; read = 0; MDRin = 0;
            end
            Reg_load3b: begin
                #10; MDRout = 1; R5in = 1;
                #15; MDRout = 0; R5in = 0;
            end
            T0: begin
                PCout = 1; MARin = 1; IncPC = 1; ZHighin = 1;
            end
            T1: begin
                Zlowout = 1; PCin = 1; read = 1; MDRin = 1;
                Mdatain <= 32'h28918000; 
            end
            T2: begin
                MDRout = 1; IRin = 1;
            end
            T3: begin
                R7out = 1; Zin = 1;
				#15 R7out = 0; Zin = 0;
            end
            T4: begin
                Zlowout = 1; R6in = 1; 
                #15 Zlowout = 0; R6in = 0; 
            end
        endcase
    end
endmodule
